library verilog;
use verilog.vl_types.all;
entity cpu_top_tb is
end cpu_top_tb;
