library verilog;
use verilog.vl_types.all;
entity reg_file_tb is
end reg_file_tb;
