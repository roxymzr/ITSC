library verilog;
use verilog.vl_types.all;
entity final_crypto_test is
end final_crypto_test;
