library verilog;
use verilog.vl_types.all;
entity professional_test is
end professional_test;
