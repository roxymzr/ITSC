library verilog;
use verilog.vl_types.all;
entity final_test is
end final_test;
